`define G_time 6'd6
`define Y_time 6'd2
`define R_time 6'd8